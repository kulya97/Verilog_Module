#File: fix_ff_loc.sv
set_property BEL DFF2 [get_cells LDCE_inst]
set_property LOC SLICE_X190Y205 [get_cells LDCE_inst]
set_property BEL CFF [get_cells FDRE_inst_ce2]
set_property LOC SLICE_X191Y205 [get_cells FDRE_inst_ce2]

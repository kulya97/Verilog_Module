//File: set_max_fanout.sv
(* MAX_FANOUT = 5 *) logic dv;
(* MAX_FANOUT = 5 *) logic [13 : 0] validForEgressFifo;

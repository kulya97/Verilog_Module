`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: NJUST
// Engineer: huangwenjie
// 
// Create Date: 2024/01/17 16:54:48
// Design Name: 
// Module Name: ISP_APB_REG_CFG
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ISP_APB_REG_CFG #(
    parameter APB_DBIT = 32,
    parameter APB_ABIT = 32,
    parameter CMD_DBIT = 8

) (
    input                                       i_clk,
    input                                       i_rstn,
    output reg                                  o_valid,
    input                                       i_ready,
    output reg [APB_DBIT+APB_ABIT+CMD_DBIT-1:0] o_data,
    output                                      o_init_done
);
  localparam CMD_WITDH = APB_DBIT + APB_ABIT + CMD_DBIT;
  localparam REG_NUM = 10;
  reg [9:0] init_reg_cnt;

  assign o_init_done = !o_valid;
  always @(posedge i_clk, negedge i_rstn) begin
    if (!i_rstn) o_valid <= 'd0;
    else if (init_reg_cnt <= REG_NUM - 1) o_valid <= 'd1;
    else o_valid <= 'd0;
  end
  /************************************************/
  //-- 握手成功发送下一个数据
  always @(posedge i_clk, negedge i_rstn) begin
    if (!i_rstn) init_reg_cnt <= 'd0;
    else if (o_valid && i_ready) init_reg_cnt <= init_reg_cnt + 1'd1;
    else init_reg_cnt <= init_reg_cnt;
  end
  //-- 表
  always @(posedge i_clk, negedge i_rstn) begin
    if (!i_rstn) begin
    end else begin
      case (init_reg_cnt)
        10'd0000: o_data <= 72'hff_0000_0001_1234_0000;
        10'd0001: o_data <= 72'hff_0000_0001_1234_0001;
        10'd0002: o_data <= 72'hff_0000_0001_1234_0002;
        10'd0003: o_data <= 72'hff_0000_0001_1234_0003;
        10'd0004: o_data <= 72'hff_0000_0001_1234_0004;
        10'd0005: o_data <= 72'hff_0000_0001_1234_0005;
        10'd0006: o_data <= 72'hff_0000_0001_1234_0006;
        10'd0007: o_data <= 72'hff_0000_0001_1234_0007;
        10'd0008: o_data <= 72'hff_0000_0001_1234_0008;
        10'd0009: o_data <= 72'hff_0000_0001_1234_0009;
        10'd0010: o_data <= 72'hff_0000_0001_1234_0010;
        10'd0011: o_data <= 72'hff_0000_0001_1234_0011;
        10'd0012: o_data <= 72'hff_0000_0001_1234_0012;
        10'd0013: o_data <= 72'hff_0000_0001_1234_0013;
        10'd0014: o_data <= 72'hff_0000_0001_1234_0014;
        10'd0015: o_data <= 72'hff_0000_0001_1234_0015;
        10'd0016: o_data <= 72'hff_0000_0001_1234_0016;
        10'd0017: o_data <= 72'hff_0000_0001_1234_0017;
        10'd0018: o_data <= 72'hff_0000_0001_1234_0018;
        10'd0019: o_data <= 72'hff_0000_0001_1234_0019;
        10'd0020: o_data <= 72'hff_0000_0001_1234_0020;
        10'd0021: o_data <= 72'hff_0000_0001_1234_0021;
        10'd0022: o_data <= 72'hff_0000_0001_1234_0022;
        10'd0023: o_data <= 72'hff_0000_0001_1234_0023;
        10'd0024: o_data <= 72'hff_0000_0001_1234_0024;
        10'd0025: o_data <= 72'hff_0000_0001_1234_0025;
        10'd0026: o_data <= 72'hff_0000_0001_1234_0026;
        10'd0027: o_data <= 72'hff_0000_0001_1234_0027;
        10'd0028: o_data <= 72'hff_0000_0001_1234_0028;
        10'd0029: o_data <= 72'hff_0000_0001_1234_0029;
        10'd0030: o_data <= 72'hff_0000_0001_1234_0030;
        10'd0031: o_data <= 72'hff_0000_0001_1234_0031;
        10'd0032: o_data <= 72'hff_0000_0001_1234_0032;
        10'd0033: o_data <= 72'hff_0000_0001_1234_0033;
        10'd0034: o_data <= 72'hff_0000_0001_1234_0034;
        10'd0035: o_data <= 72'hff_0000_0001_1234_0035;
        10'd0036: o_data <= 72'hff_0000_0001_1234_0036;
        10'd0037: o_data <= 72'hff_0000_0001_1234_0037;
        10'd0038: o_data <= 72'hff_0000_0001_1234_0038;
        10'd0039: o_data <= 72'hff_0000_0001_1234_0039;
        10'd0040: o_data <= 72'hff_0000_0001_1234_0040;
        10'd0041: o_data <= 72'hff_0000_0001_1234_0041;
        10'd0042: o_data <= 72'hff_0000_0001_1234_0042;
        10'd0043: o_data <= 72'hff_0000_0001_1234_0043;
        10'd0044: o_data <= 72'hff_0000_0001_1234_0044;
        10'd0045: o_data <= 72'hff_0000_0001_1234_0045;
        10'd0046: o_data <= 72'hff_0000_0001_1234_0046;
        10'd0047: o_data <= 72'hff_0000_0001_1234_0047;
        10'd0048: o_data <= 72'hff_0000_0001_1234_0048;
        10'd0049: o_data <= 72'hff_0000_0001_1234_0049;
        10'd0050: o_data <= 72'hff_0000_0001_1234_0050;
        10'd0051: o_data <= 72'hff_0000_0001_1234_0051;
        10'd0052: o_data <= 72'hff_0000_0001_1234_0052;
        10'd0053: o_data <= 72'hff_0000_0001_1234_0053;
        10'd0054: o_data <= 72'hff_0000_0001_1234_0054;
        10'd0055: o_data <= 72'hff_0000_0001_1234_0055;
        10'd0056: o_data <= 72'hff_0000_0001_1234_0056;
        10'd0057: o_data <= 72'hff_0000_0001_1234_0057;
        10'd0058: o_data <= 72'hff_0000_0001_1234_0058;
        10'd0059: o_data <= 72'hff_0000_0001_1234_0059;
        10'd0060: o_data <= 72'hff_0000_0001_1234_0060;
        10'd0061: o_data <= 72'hff_0000_0001_1234_0061;
        10'd0062: o_data <= 72'hff_0000_0001_1234_0062;
        10'd0063: o_data <= 72'hff_0000_0001_1234_0063;
        10'd0064: o_data <= 72'hff_0000_0001_1234_0064;
        10'd0065: o_data <= 72'hff_0000_0001_1234_0065;
        10'd0066: o_data <= 72'hff_0000_0001_1234_0066;
        10'd0067: o_data <= 72'hff_0000_0001_1234_0067;
        10'd0068: o_data <= 72'hff_0000_0001_1234_0068;
        10'd0069: o_data <= 72'hff_0000_0001_1234_0069;
        10'd0070: o_data <= 72'hff_0000_0001_1234_0070;
        10'd0071: o_data <= 72'hff_0000_0001_1234_0071;
        10'd0072: o_data <= 72'hff_0000_0001_1234_0072;
        10'd0073: o_data <= 72'hff_0000_0001_1234_0073;
        10'd0074: o_data <= 72'hff_0000_0001_1234_0074;
        10'd0075: o_data <= 72'hff_0000_0001_1234_0075;
        10'd0076: o_data <= 72'hff_0000_0001_1234_0076;
        10'd0077: o_data <= 72'hff_0000_0001_1234_0077;
        10'd0078: o_data <= 72'hff_0000_0001_1234_0078;
        10'd0079: o_data <= 72'hff_0000_0001_1234_0079;
        10'd0080: o_data <= 72'hff_0000_0001_1234_0080;
        10'd0081: o_data <= 72'hff_0000_0001_1234_0081;
        10'd0082: o_data <= 72'hff_0000_0001_1234_0082;
        10'd0083: o_data <= 72'hff_0000_0001_1234_0083;
        10'd0084: o_data <= 72'hff_0000_0001_1234_0084;
        10'd0085: o_data <= 72'hff_0000_0001_1234_0085;
        10'd0086: o_data <= 72'hff_0000_0001_1234_0086;
        10'd0087: o_data <= 72'hff_0000_0001_1234_0087;
        10'd0088: o_data <= 72'hff_0000_0001_1234_0088;
        10'd0089: o_data <= 72'hff_0000_0001_1234_0089;
        10'd0090: o_data <= 72'hff_0000_0001_1234_0090;
        10'd0091: o_data <= 72'hff_0000_0001_1234_0091;
        10'd0092: o_data <= 72'hff_0000_0001_1234_0092;
        10'd0093: o_data <= 72'hff_0000_0001_1234_0093;
        10'd0094: o_data <= 72'hff_0000_0001_1234_0094;
        10'd0095: o_data <= 72'hff_0000_0001_1234_0095;
        10'd0096: o_data <= 72'hff_0000_0001_1234_0096;
        10'd0097: o_data <= 72'hff_0000_0001_1234_0097;
        10'd0098: o_data <= 72'hff_0000_0001_1234_0098;
        10'd0099: o_data <= 72'hff_0000_0001_1234_0099;
        10'd0100: o_data <= 72'hff_0000_0001_1234_0100;
        10'd0101: o_data <= 72'hff_0000_0001_1234_0101;
        10'd0102: o_data <= 72'hff_0000_0001_1234_0102;
        10'd0103: o_data <= 72'hff_0000_0001_1234_0103;
        10'd0104: o_data <= 72'hff_0000_0001_1234_0104;
        10'd0105: o_data <= 72'hff_0000_0001_1234_0105;
        10'd0106: o_data <= 72'hff_0000_0001_1234_0106;
        10'd0107: o_data <= 72'hff_0000_0001_1234_0107;
        10'd0108: o_data <= 72'hff_0000_0001_1234_0108;
        10'd0109: o_data <= 72'hff_0000_0001_1234_0109;
        10'd0110: o_data <= 72'hff_0000_0001_1234_0110;
        10'd0111: o_data <= 72'hff_0000_0001_1234_0111;
        10'd0112: o_data <= 72'hff_0000_0001_1234_0112;
        10'd0113: o_data <= 72'hff_0000_0001_1234_0113;
        10'd0114: o_data <= 72'hff_0000_0001_1234_0114;
        10'd0115: o_data <= 72'hff_0000_0001_1234_0115;
        10'd0116: o_data <= 72'hff_0000_0001_1234_0116;
        10'd0117: o_data <= 72'hff_0000_0001_1234_0117;
        10'd0118: o_data <= 72'hff_0000_0001_1234_0118;
        10'd0119: o_data <= 72'hff_0000_0001_1234_0119;
        10'd0120: o_data <= 72'hff_0000_0001_1234_0120;
        10'd0121: o_data <= 72'hff_0000_0001_1234_0121;
        10'd0122: o_data <= 72'hff_0000_0001_1234_0122;
        10'd0123: o_data <= 72'hff_0000_0001_1234_0123;
        10'd0124: o_data <= 72'hff_0000_0001_1234_0124;
        10'd0125: o_data <= 72'hff_0000_0001_1234_0125;
        10'd0126: o_data <= 72'hff_0000_0001_1234_0126;
        10'd0127: o_data <= 72'hff_0000_0001_1234_0127;
        10'd0128: o_data <= 72'hff_0000_0001_1234_0128;
        10'd0129: o_data <= 72'hff_0000_0001_1234_0129;
        10'd0130: o_data <= 72'hff_0000_0001_1234_0130;
        10'd0131: o_data <= 72'hff_0000_0001_1234_0131;
        10'd0132: o_data <= 72'hff_0000_0001_1234_0132;
        10'd0133: o_data <= 72'hff_0000_0001_1234_0133;
        10'd0134: o_data <= 72'hff_0000_0001_1234_0134;
        10'd0135: o_data <= 72'hff_0000_0001_1234_0135;
        10'd0136: o_data <= 72'hff_0000_0001_1234_0136;
        10'd0137: o_data <= 72'hff_0000_0001_1234_0137;
        10'd0138: o_data <= 72'hff_0000_0001_1234_0138;
        10'd0139: o_data <= 72'hff_0000_0001_1234_0139;
        10'd0140: o_data <= 72'hff_0000_0001_1234_0140;
        10'd0141: o_data <= 72'hff_0000_0001_1234_0141;
        10'd0142: o_data <= 72'hff_0000_0001_1234_0142;
        10'd0143: o_data <= 72'hff_0000_0001_1234_0143;
        10'd0144: o_data <= 72'hff_0000_0001_1234_0144;
        10'd0145: o_data <= 72'hff_0000_0001_1234_0145;
        10'd0146: o_data <= 72'hff_0000_0001_1234_0146;
        10'd0147: o_data <= 72'hff_0000_0001_1234_0147;
        10'd0148: o_data <= 72'hff_0000_0001_1234_0148;
        10'd0149: o_data <= 72'hff_0000_0001_1234_0149;
        10'd0150: o_data <= 72'hff_0000_0001_1234_0150;
        10'd0151: o_data <= 72'hff_0000_0001_1234_0151;
        10'd0152: o_data <= 72'hff_0000_0001_1234_0152;
        10'd0153: o_data <= 72'hff_0000_0001_1234_0153;
        10'd0154: o_data <= 72'hff_0000_0001_1234_0154;
        10'd0155: o_data <= 72'hff_0000_0001_1234_0155;
        10'd0156: o_data <= 72'hff_0000_0001_1234_0156;
        10'd0157: o_data <= 72'hff_0000_0001_1234_0157;
        10'd0158: o_data <= 72'hff_0000_0001_1234_0158;
        10'd0159: o_data <= 72'hff_0000_0001_1234_0159;
        10'd0160: o_data <= 72'hff_0000_0001_1234_0160;
        10'd0161: o_data <= 72'hff_0000_0001_1234_0161;
        10'd0162: o_data <= 72'hff_0000_0001_1234_0162;
        10'd0163: o_data <= 72'hff_0000_0001_1234_0163;
        10'd0164: o_data <= 72'hff_0000_0001_1234_0164;
        10'd0165: o_data <= 72'hff_0000_0001_1234_0165;
        10'd0166: o_data <= 72'hff_0000_0001_1234_0166;
        10'd0167: o_data <= 72'hff_0000_0001_1234_0167;
        10'd0168: o_data <= 72'hff_0000_0001_1234_0168;
        10'd0169: o_data <= 72'hff_0000_0001_1234_0169;
        10'd0170: o_data <= 72'hff_0000_0001_1234_0170;
        10'd0171: o_data <= 72'hff_0000_0001_1234_0171;
        10'd0172: o_data <= 72'hff_0000_0001_1234_0172;
        10'd0173: o_data <= 72'hff_0000_0001_1234_0173;
        10'd0174: o_data <= 72'hff_0000_0001_1234_0174;
        10'd0175: o_data <= 72'hff_0000_0001_1234_0175;
        10'd0176: o_data <= 72'hff_0000_0001_1234_0176;
        10'd0177: o_data <= 72'hff_0000_0001_1234_0177;
        10'd0178: o_data <= 72'hff_0000_0001_1234_0178;
        10'd0179: o_data <= 72'hff_0000_0001_1234_0179;
        10'd0180: o_data <= 72'hff_0000_0001_1234_0180;
        10'd0181: o_data <= 72'hff_0000_0001_1234_0181;
        10'd0182: o_data <= 72'hff_0000_0001_1234_0182;
        10'd0183: o_data <= 72'hff_0000_0001_1234_0183;
        10'd0184: o_data <= 72'hff_0000_0001_1234_0184;
        10'd0185: o_data <= 72'hff_0000_0001_1234_0185;
        10'd0186: o_data <= 72'hff_0000_0001_1234_0186;
        10'd0187: o_data <= 72'hff_0000_0001_1234_0187;
        10'd0188: o_data <= 72'hff_0000_0001_1234_0188;
        10'd0189: o_data <= 72'hff_0000_0001_1234_0189;
        10'd0190: o_data <= 72'hff_0000_0001_1234_0190;
        10'd0191: o_data <= 72'hff_0000_0001_1234_0191;
        10'd0192: o_data <= 72'hff_0000_0001_1234_0192;
        10'd0193: o_data <= 72'hff_0000_0001_1234_0193;
        10'd0194: o_data <= 72'hff_0000_0001_1234_0194;
        10'd0195: o_data <= 72'hff_0000_0001_1234_0195;
        10'd0196: o_data <= 72'hff_0000_0001_1234_0196;
        10'd0197: o_data <= 72'hff_0000_0001_1234_0197;
        10'd0198: o_data <= 72'hff_0000_0001_1234_0198;
        10'd0199: o_data <= 72'hff_0000_0001_1234_0199;
        10'd0200: o_data <= 72'hff_0000_0001_1234_0200;
        10'd0201: o_data <= 72'hff_0000_0001_1234_0201;
        10'd0202: o_data <= 72'hff_0000_0001_1234_0202;
        10'd0203: o_data <= 72'hff_0000_0001_1234_0203;
        10'd0204: o_data <= 72'hff_0000_0001_1234_0204;
        10'd0205: o_data <= 72'hff_0000_0001_1234_0205;
        10'd0206: o_data <= 72'hff_0000_0001_1234_0206;
        10'd0207: o_data <= 72'hff_0000_0001_1234_0207;
        10'd0208: o_data <= 72'hff_0000_0001_1234_0208;
        10'd0209: o_data <= 72'hff_0000_0001_1234_0209;
        10'd0210: o_data <= 72'hff_0000_0001_1234_0210;
        10'd0211: o_data <= 72'hff_0000_0001_1234_0211;
        10'd0212: o_data <= 72'hff_0000_0001_1234_0212;
        10'd0213: o_data <= 72'hff_0000_0001_1234_0213;
        10'd0214: o_data <= 72'hff_0000_0001_1234_0214;
        10'd0215: o_data <= 72'hff_0000_0001_1234_0215;
        10'd0216: o_data <= 72'hff_0000_0001_1234_0216;
        10'd0217: o_data <= 72'hff_0000_0001_1234_0217;
        10'd0218: o_data <= 72'hff_0000_0001_1234_0218;
        10'd0219: o_data <= 72'hff_0000_0001_1234_0219;
        10'd0220: o_data <= 72'hff_0000_0001_1234_0220;
        10'd0221: o_data <= 72'hff_0000_0001_1234_0221;
        10'd0222: o_data <= 72'hff_0000_0001_1234_0222;
        10'd0223: o_data <= 72'hff_0000_0001_1234_0223;
        10'd0224: o_data <= 72'hff_0000_0001_1234_0224;
        10'd0225: o_data <= 72'hff_0000_0001_1234_0225;
        10'd0226: o_data <= 72'hff_0000_0001_1234_0226;
        10'd0227: o_data <= 72'hff_0000_0001_1234_0227;
        10'd0228: o_data <= 72'hff_0000_0001_1234_0228;
        10'd0229: o_data <= 72'hff_0000_0001_1234_0229;
        10'd0230: o_data <= 72'hff_0000_0001_1234_0230;
        10'd0231: o_data <= 72'hff_0000_0001_1234_0231;
        10'd0232: o_data <= 72'hff_0000_0001_1234_0232;
        10'd0233: o_data <= 72'hff_0000_0001_1234_0233;
        10'd0234: o_data <= 72'hff_0000_0001_1234_0234;
        10'd0235: o_data <= 72'hff_0000_0001_1234_0235;
        10'd0236: o_data <= 72'hff_0000_0001_1234_0236;
        10'd0237: o_data <= 72'hff_0000_0001_1234_0237;
        10'd0238: o_data <= 72'hff_0000_0001_1234_0238;
        10'd0239: o_data <= 72'hff_0000_0001_1234_0239;
        10'd0240: o_data <= 72'hff_0000_0001_1234_0240;
        10'd0241: o_data <= 72'hff_0000_0001_1234_0241;
        10'd0242: o_data <= 72'hff_0000_0001_1234_0242;
        10'd0243: o_data <= 72'hff_0000_0001_1234_0243;
        10'd0244: o_data <= 72'hff_0000_0001_1234_0244;
        10'd0245: o_data <= 72'hff_0000_0001_1234_0245;
        10'd0246: o_data <= 72'hff_0000_0001_1234_0246;
        10'd0247: o_data <= 72'hff_0000_0001_1234_0247;
        10'd0248: o_data <= 72'hff_0000_0001_1234_0248;
        10'd0249: o_data <= 72'hff_0000_0001_1234_0249;
        10'd0250: o_data <= 72'hff_0000_0001_1234_0250;
        10'd0251: o_data <= 72'hff_0000_0001_1234_0251;
        10'd0252: o_data <= 72'hff_0000_0001_1234_0252;
        10'd0253: o_data <= 72'hff_0000_0001_1234_0253;
        10'd0254: o_data <= 72'hff_0000_0001_1234_0254;
        default:  o_data <= 72'hff_0000_0001_1234_0254;
      endcase
    end
  end
endmodule
